library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity g89_FSM is 
	
	Port (
		enable		: in	std_logic;			-- FSM will only work if enable is 1
		direction 	: in	std_logic;			-- FSM will go with 2 directions {'0': right, '1': left}
		reset		: in  	std_logic;			-- FSM will be reset if reset is 0
		clk		: in 	std_logic;			-- FSM will only be active when at the rising edge of the clk
		count		: out 	std_logic_vector (3 downto 0)	-- This represents the current state of the FSM
	);
	
end g89_FSM;

architecture behaviour of g89_FSM is

	type State_type 	is	(A, B, C, D, E, F, G, H, I, J, K, L, M, N, O);
	signal present_state	: 	State_type;
	signal temp		:	std_logic_vector (3 downto 0);

begin 
	process(enable, direction, reset, clk)
	begin 
	
	if (reset = '0') then 					-- Reset FSM when reset is 0
		present_state <= A;
			
	elsif (rising_edge(clk) and enable = '1') then		-- FSM opreates at the rising edge of clk and when enable is 1
		case present_state is 
			when A => 
				if direction = '0' then	
					present_state <= B;
				else 
					present_state <= O;
				end if;
						
			when B => 
				if direction = '0' then 
					present_state <= C;
				else 
					present_state <= A;
				end if;
						
			when C => 
				if direction = '0' then
					present_state <= D;
				else 
					present_state <= B;
				end if;
						
			when D => 
				if direction = '0' then
					present_state <= E;
				else 
					present_state <= C;
				end if;
						
			when E => 
				if direction = '0' then
					present_state <= F;
				else 
					present_state <= D;
				end if;
						
			when F => 
				if direction = '0' then
					present_state <= G;
				else 
					present_state <= E;
				end if;
					
			when G => 
				if direction = '0' then
					present_state <= H;
				else 
					present_state <= F;
				end if;
						
			when H => 
				if direction = '0' then
					present_state <= I;
				else 
					present_state <= G;
				end if;
					
			when I => 
				if direction = '0' then
					present_state <= J;
				else 
					present_state <= H;
				end if;
						
			when J => 
				if direction = '0' then
					present_state <= K;
				else 
					present_state <= I;
				end if;
					
			when K => 
				if direction = '0' then
					present_state <= L;
				else 
					present_state <= J;
				end if;
						
			when L => 
				if direction = '0' then
					present_state <= M;
				else 
					present_state <= K;
				end if;
					
			when M => 
				if direction = '0' then
					present_state <= N;
				else 
					present_state <= L;
				end if;
						
			when N => 
				if direction = '0' then
					present_state <= O;
				else 
					present_state <= M;
				end if;
						
			when O => 
				if direction = '0' then
					present_state <= A;
				else 
					present_state <= N;
				end if;
			end case;
			
	end if;
	
	case present_state is 
		when A => temp <= "0001";
		when B => temp <= "0010";
		when C => temp <= "0100";
		when D => temp <= "1000";
		when E => temp <= "0011";
		when F => temp <= "0110";
		when G => temp <= "1100";
		when H => temp <= "1011";
		when I => temp <= "0101";
		when J => temp <= "1010";
		when K => temp <= "0111";
		when L => temp <= "1110";
		when M => temp <= "1111";
		when N => temp <= "1101";
		when O => temp <= "1001";
		when others => temp <= "0000";
	end case;
			
	end process;
	count <= temp;
end behaviour;
		
			
			
			
			
			
			
			
			
							
